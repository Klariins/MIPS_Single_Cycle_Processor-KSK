module InstructionMemory (read_Address, instruction, clock);

	input [31:0] read_Address;
	input clock;
	output [31:0] instruction;
	reg [75:0] Memory [75:0];
	integer flag_Start = 1;
	
	always@(posedge clock)
	begin
		if (flag_Start == 1)
		begin	
		
			Memory[0] = 32'b100110_00000_00001_0000000000000000;		// in r[1]
			Memory[1] = 32'b011110_00000_00001_0000000000000001;		// Mem[1] = r[1]
			Memory[2] = 32'b100111_00000000000000000000000001;			// out d[1]
			Memory[3] = 32'b100110_00000_00010_0000000000000000;		// in r[2]
			Memory[4] = 32'b011110_00000_00010_0000000000000010;		// Mem[2] = r[2]
			Memory[5] = 32'b100111_00000000000000000000000010;			// out d[2]
			Memory[6] = 32'b000001_00011_00011_0000000000000001;		// r[3] = r[3] + 1 (r[3] = Im(1))
			Memory[7] = 32'b100010_00000000000000000000011110;			// jal 30
			Memory[8] = 32'b011101_00000_00100_0000000000000001;		// r[4] = Mem[1] 100000_00001_00100_0000000000000000;
			Memory[9] = 32'b000100_00100_00001_00100_00000000000;		// r[4] = r[4] * r[1]
			Memory[10] = 32'b000010_00010_00011_00010_00000000000; 	// r[2] = r[2] - r[3]
			Memory[11] = 32'b010100_00010_00011_0000000000001001; 	// r[2] > r[3], PC = 9
			Memory[12] = 32'b100001_00000000000000000000111100;		// j 60
			
			Memory[30] = 32'b010000_00000_00010_0000000000101000; 	// r[2] == r[0], PC = 40 
			Memory[31] = 32'b010000_00010_00011_0000000000110010; 	// r[2] == r[3], PC = 50
			Memory[32] = 32'b100011_11111_000000000000000000000;		// jr 31
			
			Memory[40] = 32'b011110_00000_00011_0000000000000011;		// Mem[3] = r[3]
			Memory[41] = 32'b100111_00000000000000000000000011;		// out d[3]
			Memory[42] = 32'b100001_00000000000000000001000110;		// j 70
			
			Memory[50] = 32'b011110_00000_00001_0000000000000011;		// Mem[3] = r[1]
			Memory[51] = 32'b100111_00000000000000000000000011;		// out d[3]
			Memory[52] = 32'b100001_00000000000000000001000110;		// j 70
			
			Memory[60] = 32'b011110_00000_00100_0000000000000100;		// Mem[4] = r[4]
			Memory[61] = 32'b100111_00000000000000000000000100;		// out d[4]
			Memory[62] = 32'b100001_00000000000000000001000110;		// j 70
			
			Memory[70] = 32'b100101_00000000000000000000000000;    	// halt
 
			flag_Start <= 0;
		end
	end
	
	assign instruction = Memory[read_Address];	
	
endmodule
